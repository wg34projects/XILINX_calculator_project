--
-- FHTW - BEL3 - DSD - calculator project
--
--
-- Author:	Helmut Resch
--			el16b005
--			BEL3
--
-- File:	tb_io_ctrl_.vhd
--
-- Version history:
--
-- v_0.1	13.11.2017	IO Ctrl + Testbench
-- v_0.2	15.11.2017	Calc Ctrl + Testbench
--
-- Design Unit:	IO Control Unit Testbench
--				Entity
--
-- Description:	The IO Control unit is part of the calculator project.
--				It manages the interface to the 7-segment displays,
--				the LEDs, the push buttons and the switches of the
--				Digilent Basys3 FPGA board.
--
--
-- below doxygen documentation blocks

--! @file tb_io_ctrl_.vhd
--! @brief IO Control Unit Testbench Entity

library IEEE;
use IEEE.std_logic_1164.all;

--! @brief IO Control Unit Testbench Entity
--! @details The IO Control unit is part of the calculator project.

entity tb_io_ctrl is

end tb_io_ctrl;
